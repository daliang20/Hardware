// sys_vga.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module sys_vga (
		input  wire        alt_vip_itc_0_clocked_video_vid_clk,       // alt_vip_itc_0_clocked_video.vid_clk
		output wire [31:0] alt_vip_itc_0_clocked_video_vid_data,      //                            .vid_data
		output wire        alt_vip_itc_0_clocked_video_underflow,     //                            .underflow
		output wire        alt_vip_itc_0_clocked_video_vid_datavalid, //                            .vid_datavalid
		output wire        alt_vip_itc_0_clocked_video_vid_v_sync,    //                            .vid_v_sync
		output wire        alt_vip_itc_0_clocked_video_vid_h_sync,    //                            .vid_h_sync
		output wire        alt_vip_itc_0_clocked_video_vid_f,         //                            .vid_f
		output wire        alt_vip_itc_0_clocked_video_vid_h,         //                            .vid_h
		output wire        alt_vip_itc_0_clocked_video_vid_v,         //                            .vid_v
		output wire        clk_65_clk,                                //                      clk_65.clk
		input  wire        clock_bridge_0_in_clk_clk,                 //       clock_bridge_0_in_clk.clk
		input  wire [31:0] fifo_fpga_to_hps_in_writedata,             //         fifo_fpga_to_hps_in.writedata
		input  wire        fifo_fpga_to_hps_in_write,                 //                            .write
		output wire        fifo_fpga_to_hps_in_waitrequest,           //                            .waitrequest
		input  wire [2:0]  fifo_fpga_to_hps_in_csr_address,           //     fifo_fpga_to_hps_in_csr.address
		input  wire        fifo_fpga_to_hps_in_csr_read,              //                            .read
		input  wire [31:0] fifo_fpga_to_hps_in_csr_writedata,         //                            .writedata
		input  wire        fifo_fpga_to_hps_in_csr_write,             //                            .write
		output wire [31:0] fifo_fpga_to_hps_in_csr_readdata,          //                            .readdata
		output wire [31:0] fifo_hps_to_fpga_out_readdata,             //        fifo_hps_to_fpga_out.readdata
		input  wire        fifo_hps_to_fpga_out_read,                 //                            .read
		output wire        fifo_hps_to_fpga_out_waitrequest,          //                            .waitrequest
		input  wire [2:0]  fifo_hps_to_fpga_out_csr_address,          //    fifo_hps_to_fpga_out_csr.address
		input  wire        fifo_hps_to_fpga_out_csr_read,             //                            .read
		input  wire [31:0] fifo_hps_to_fpga_out_csr_writedata,        //                            .writedata
		input  wire        fifo_hps_to_fpga_out_csr_write,            //                            .write
		output wire [31:0] fifo_hps_to_fpga_out_csr_readdata,         //                            .readdata
		output wire [31:0] hex5_0bus_export,                          //                   hex5_0bus.export
		inout  wire        hps_io_hps_io_sdio_inst_CMD,               //                      hps_io.hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,                //                            .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,                //                            .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,               //                            .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,                //                            .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,                //                            .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,                //                            .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,                //                            .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,                //                            .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,                //                            .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,                //                            .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,                //                            .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,                //                            .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,                //                            .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,               //                            .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,               //                            .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,               //                            .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,               //                            .hps_io_usb1_inst_NXT
		input  wire        hps_io_hps_io_uart0_inst_RX,               //                            .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,               //                            .hps_io_uart0_inst_TX
		output wire [14:0] memory_mem_a,                              //                      memory.mem_a
		output wire [2:0]  memory_mem_ba,                             //                            .mem_ba
		output wire        memory_mem_ck,                             //                            .mem_ck
		output wire        memory_mem_ck_n,                           //                            .mem_ck_n
		output wire        memory_mem_cke,                            //                            .mem_cke
		output wire        memory_mem_cs_n,                           //                            .mem_cs_n
		output wire        memory_mem_ras_n,                          //                            .mem_ras_n
		output wire        memory_mem_cas_n,                          //                            .mem_cas_n
		output wire        memory_mem_we_n,                           //                            .mem_we_n
		output wire        memory_mem_reset_n,                        //                            .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                             //                            .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                            //                            .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                          //                            .mem_dqs_n
		output wire        memory_mem_odt,                            //                            .mem_odt
		output wire [3:0]  memory_mem_dm,                             //                            .mem_dm
		input  wire        memory_oct_rzqin,                          //                            .oct_rzqin
		input  wire [3:0]  pushbutton_export,                         //                  pushbutton.export
		input  wire [10:0] ram_s2_address,                            //                      ram_s2.address
		input  wire        ram_s2_chipselect,                         //                            .chipselect
		input  wire        ram_s2_clken,                              //                            .clken
		input  wire        ram_s2_write,                              //                            .write
		output wire [31:0] ram_s2_readdata,                           //                            .readdata
		input  wire [31:0] ram_s2_writedata,                          //                            .writedata
		input  wire [3:0]  ram_s2_byteenable,                         //                            .byteenable
		output wire        sdram_clk_clk,                             //                   sdram_clk.clk
		output wire [12:0] sdram_wire_addr,                           //                  sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                             //                            .ba
		output wire        sdram_wire_cas_n,                          //                            .cas_n
		output wire        sdram_wire_cke,                            //                            .cke
		output wire        sdram_wire_cs_n,                           //                            .cs_n
		inout  wire [15:0] sdram_wire_dq,                             //                            .dq
		output wire [1:0]  sdram_wire_dqm,                            //                            .dqm
		output wire        sdram_wire_ras_n,                          //                            .ras_n
		output wire        sdram_wire_we_n,                           //                            .we_n
		input  wire        system_ref_clk_clk,                        //              system_ref_clk.clk
		input  wire        system_ref_reset_reset,                    //            system_ref_reset.reset
		output wire [31:0] to_hex_to_led_readdata                     //               to_hex_to_led.readdata
	);

	wire          alt_vip_vfr_0_avalon_streaming_source_valid;                          // alt_vip_vfr_0:dout_valid -> alt_vip_itc_0:is_valid
	wire   [31:0] alt_vip_vfr_0_avalon_streaming_source_data;                           // alt_vip_vfr_0:dout_data -> alt_vip_itc_0:is_data
	wire          alt_vip_vfr_0_avalon_streaming_source_ready;                          // alt_vip_itc_0:is_ready -> alt_vip_vfr_0:dout_ready
	wire          alt_vip_vfr_0_avalon_streaming_source_startofpacket;                  // alt_vip_vfr_0:dout_startofpacket -> alt_vip_itc_0:is_sop
	wire          alt_vip_vfr_0_avalon_streaming_source_endofpacket;                    // alt_vip_vfr_0:dout_endofpacket -> alt_vip_itc_0:is_eop
	wire          pll_0_outclk0_clk;                                                    // pll_0:outclk_0 -> [alt_vip_itc_0:is_clk, alt_vip_vfr_0:clock, mm_interconnect_2:pll_0_outclk0_clk, rst_controller:clk]
	wire          sys_sdram_pll_0_sys_clk_clk;                                          // sys_sdram_pll_0:sys_clk_clk -> [Arm_A9_HPS:f2h_axi_clk, Arm_A9_HPS:h2f_axi_clk, Arm_A9_HPS:h2f_lw_axi_clk, alt_vip_vfr_0:master_clock, fifo_fpga_to_hps:rdclock, fifo_hps_to_fpga:wrclock, hex5_hex0:clk, mm_interconnect_0:sys_sdram_pll_0_sys_clk_clk, mm_interconnect_1:sys_sdram_pll_0_sys_clk_clk, mm_interconnect_2:sys_sdram_pll_0_sys_clk_clk, new_sdram_controller_0:clk, pll_0:refclk, pll_1:refclk, pushbuttons:clk, ram:clk, reg32_avalon_interface_0:clk, rst_controller_001:clk, rst_controller_003:clk, rst_controller_004:clk, sysid_qsys_0:clock, system_console:clk]
	wire          sys_sdram_pll_0_reset_source_reset;                                   // sys_sdram_pll_0:reset_source_reset -> [pll_0:rst, pll_1:rst, rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in1, rst_controller_003:reset_in1]
	wire  [127:0] alt_vip_vfr_0_avalon_master_readdata;                                 // mm_interconnect_0:alt_vip_vfr_0_avalon_master_readdata -> alt_vip_vfr_0:master_readdata
	wire          alt_vip_vfr_0_avalon_master_waitrequest;                              // mm_interconnect_0:alt_vip_vfr_0_avalon_master_waitrequest -> alt_vip_vfr_0:master_waitrequest
	wire   [31:0] alt_vip_vfr_0_avalon_master_address;                                  // alt_vip_vfr_0:master_address -> mm_interconnect_0:alt_vip_vfr_0_avalon_master_address
	wire          alt_vip_vfr_0_avalon_master_read;                                     // alt_vip_vfr_0:master_read -> mm_interconnect_0:alt_vip_vfr_0_avalon_master_read
	wire          alt_vip_vfr_0_avalon_master_readdatavalid;                            // mm_interconnect_0:alt_vip_vfr_0_avalon_master_readdatavalid -> alt_vip_vfr_0:master_readdatavalid
	wire    [5:0] alt_vip_vfr_0_avalon_master_burstcount;                               // alt_vip_vfr_0:master_burstcount -> mm_interconnect_0:alt_vip_vfr_0_avalon_master_burstcount
	wire    [1:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awburst;                   // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_awburst -> Arm_A9_HPS:f2h_AWBURST
	wire    [4:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awuser;                    // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_awuser -> Arm_A9_HPS:f2h_AWUSER
	wire    [3:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arlen;                     // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_arlen -> Arm_A9_HPS:f2h_ARLEN
	wire    [7:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wstrb;                     // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_wstrb -> Arm_A9_HPS:f2h_WSTRB
	wire          mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wready;                    // Arm_A9_HPS:f2h_WREADY -> mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_wready
	wire    [7:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rid;                       // Arm_A9_HPS:f2h_RID -> mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_rid
	wire          mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rready;                    // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_rready -> Arm_A9_HPS:f2h_RREADY
	wire    [3:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awlen;                     // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_awlen -> Arm_A9_HPS:f2h_AWLEN
	wire    [7:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wid;                       // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_wid -> Arm_A9_HPS:f2h_WID
	wire    [3:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arcache;                   // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_arcache -> Arm_A9_HPS:f2h_ARCACHE
	wire          mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wvalid;                    // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_wvalid -> Arm_A9_HPS:f2h_WVALID
	wire   [31:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_araddr;                    // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_araddr -> Arm_A9_HPS:f2h_ARADDR
	wire    [2:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arprot;                    // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_arprot -> Arm_A9_HPS:f2h_ARPROT
	wire    [2:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awprot;                    // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_awprot -> Arm_A9_HPS:f2h_AWPROT
	wire   [63:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wdata;                     // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_wdata -> Arm_A9_HPS:f2h_WDATA
	wire          mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arvalid;                   // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_arvalid -> Arm_A9_HPS:f2h_ARVALID
	wire    [3:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awcache;                   // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_awcache -> Arm_A9_HPS:f2h_AWCACHE
	wire    [7:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arid;                      // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_arid -> Arm_A9_HPS:f2h_ARID
	wire    [1:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arlock;                    // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_arlock -> Arm_A9_HPS:f2h_ARLOCK
	wire    [1:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awlock;                    // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_awlock -> Arm_A9_HPS:f2h_AWLOCK
	wire   [31:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awaddr;                    // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_awaddr -> Arm_A9_HPS:f2h_AWADDR
	wire    [1:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bresp;                     // Arm_A9_HPS:f2h_BRESP -> mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_bresp
	wire          mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arready;                   // Arm_A9_HPS:f2h_ARREADY -> mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_arready
	wire   [63:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rdata;                     // Arm_A9_HPS:f2h_RDATA -> mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_rdata
	wire          mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awready;                   // Arm_A9_HPS:f2h_AWREADY -> mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_awready
	wire    [1:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arburst;                   // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_arburst -> Arm_A9_HPS:f2h_ARBURST
	wire    [2:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arsize;                    // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_arsize -> Arm_A9_HPS:f2h_ARSIZE
	wire          mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bready;                    // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_bready -> Arm_A9_HPS:f2h_BREADY
	wire          mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rlast;                     // Arm_A9_HPS:f2h_RLAST -> mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_rlast
	wire          mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wlast;                     // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_wlast -> Arm_A9_HPS:f2h_WLAST
	wire    [1:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rresp;                     // Arm_A9_HPS:f2h_RRESP -> mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_rresp
	wire    [7:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awid;                      // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_awid -> Arm_A9_HPS:f2h_AWID
	wire    [7:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bid;                       // Arm_A9_HPS:f2h_BID -> mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_bid
	wire          mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bvalid;                    // Arm_A9_HPS:f2h_BVALID -> mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_bvalid
	wire    [2:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awsize;                    // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_awsize -> Arm_A9_HPS:f2h_AWSIZE
	wire          mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awvalid;                   // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_awvalid -> Arm_A9_HPS:f2h_AWVALID
	wire    [4:0] mm_interconnect_0_arm_a9_hps_f2h_axi_slave_aruser;                    // mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_aruser -> Arm_A9_HPS:f2h_ARUSER
	wire          mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rvalid;                    // Arm_A9_HPS:f2h_RVALID -> mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_rvalid
	wire    [1:0] arm_a9_hps_h2f_axi_master_awburst;                                    // Arm_A9_HPS:h2f_AWBURST -> mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_awburst
	wire    [3:0] arm_a9_hps_h2f_axi_master_arlen;                                      // Arm_A9_HPS:h2f_ARLEN -> mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_arlen
	wire   [15:0] arm_a9_hps_h2f_axi_master_wstrb;                                      // Arm_A9_HPS:h2f_WSTRB -> mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_wstrb
	wire          arm_a9_hps_h2f_axi_master_wready;                                     // mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_wready -> Arm_A9_HPS:h2f_WREADY
	wire   [11:0] arm_a9_hps_h2f_axi_master_rid;                                        // mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_rid -> Arm_A9_HPS:h2f_RID
	wire          arm_a9_hps_h2f_axi_master_rready;                                     // Arm_A9_HPS:h2f_RREADY -> mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_rready
	wire    [3:0] arm_a9_hps_h2f_axi_master_awlen;                                      // Arm_A9_HPS:h2f_AWLEN -> mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_awlen
	wire   [11:0] arm_a9_hps_h2f_axi_master_wid;                                        // Arm_A9_HPS:h2f_WID -> mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_wid
	wire    [3:0] arm_a9_hps_h2f_axi_master_arcache;                                    // Arm_A9_HPS:h2f_ARCACHE -> mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_arcache
	wire          arm_a9_hps_h2f_axi_master_wvalid;                                     // Arm_A9_HPS:h2f_WVALID -> mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_wvalid
	wire   [29:0] arm_a9_hps_h2f_axi_master_araddr;                                     // Arm_A9_HPS:h2f_ARADDR -> mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_araddr
	wire    [2:0] arm_a9_hps_h2f_axi_master_arprot;                                     // Arm_A9_HPS:h2f_ARPROT -> mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_arprot
	wire    [2:0] arm_a9_hps_h2f_axi_master_awprot;                                     // Arm_A9_HPS:h2f_AWPROT -> mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_awprot
	wire  [127:0] arm_a9_hps_h2f_axi_master_wdata;                                      // Arm_A9_HPS:h2f_WDATA -> mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_wdata
	wire          arm_a9_hps_h2f_axi_master_arvalid;                                    // Arm_A9_HPS:h2f_ARVALID -> mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_arvalid
	wire    [3:0] arm_a9_hps_h2f_axi_master_awcache;                                    // Arm_A9_HPS:h2f_AWCACHE -> mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_awcache
	wire   [11:0] arm_a9_hps_h2f_axi_master_arid;                                       // Arm_A9_HPS:h2f_ARID -> mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_arid
	wire    [1:0] arm_a9_hps_h2f_axi_master_arlock;                                     // Arm_A9_HPS:h2f_ARLOCK -> mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_arlock
	wire    [1:0] arm_a9_hps_h2f_axi_master_awlock;                                     // Arm_A9_HPS:h2f_AWLOCK -> mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_awlock
	wire   [29:0] arm_a9_hps_h2f_axi_master_awaddr;                                     // Arm_A9_HPS:h2f_AWADDR -> mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_awaddr
	wire    [1:0] arm_a9_hps_h2f_axi_master_bresp;                                      // mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_bresp -> Arm_A9_HPS:h2f_BRESP
	wire          arm_a9_hps_h2f_axi_master_arready;                                    // mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_arready -> Arm_A9_HPS:h2f_ARREADY
	wire  [127:0] arm_a9_hps_h2f_axi_master_rdata;                                      // mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_rdata -> Arm_A9_HPS:h2f_RDATA
	wire          arm_a9_hps_h2f_axi_master_awready;                                    // mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_awready -> Arm_A9_HPS:h2f_AWREADY
	wire    [1:0] arm_a9_hps_h2f_axi_master_arburst;                                    // Arm_A9_HPS:h2f_ARBURST -> mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_arburst
	wire    [2:0] arm_a9_hps_h2f_axi_master_arsize;                                     // Arm_A9_HPS:h2f_ARSIZE -> mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_arsize
	wire          arm_a9_hps_h2f_axi_master_bready;                                     // Arm_A9_HPS:h2f_BREADY -> mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_bready
	wire          arm_a9_hps_h2f_axi_master_rlast;                                      // mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_rlast -> Arm_A9_HPS:h2f_RLAST
	wire          arm_a9_hps_h2f_axi_master_wlast;                                      // Arm_A9_HPS:h2f_WLAST -> mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_wlast
	wire    [1:0] arm_a9_hps_h2f_axi_master_rresp;                                      // mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_rresp -> Arm_A9_HPS:h2f_RRESP
	wire   [11:0] arm_a9_hps_h2f_axi_master_awid;                                       // Arm_A9_HPS:h2f_AWID -> mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_awid
	wire   [11:0] arm_a9_hps_h2f_axi_master_bid;                                        // mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_bid -> Arm_A9_HPS:h2f_BID
	wire          arm_a9_hps_h2f_axi_master_bvalid;                                     // mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_bvalid -> Arm_A9_HPS:h2f_BVALID
	wire    [2:0] arm_a9_hps_h2f_axi_master_awsize;                                     // Arm_A9_HPS:h2f_AWSIZE -> mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_awsize
	wire          arm_a9_hps_h2f_axi_master_awvalid;                                    // Arm_A9_HPS:h2f_AWVALID -> mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_awvalid
	wire          arm_a9_hps_h2f_axi_master_rvalid;                                     // mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_rvalid -> Arm_A9_HPS:h2f_RVALID
	wire          mm_interconnect_1_fifo_hps_to_fpga_in_waitrequest;                    // fifo_hps_to_fpga:avalonmm_write_slave_waitrequest -> mm_interconnect_1:fifo_hps_to_fpga_in_waitrequest
	wire          mm_interconnect_1_fifo_hps_to_fpga_in_write;                          // mm_interconnect_1:fifo_hps_to_fpga_in_write -> fifo_hps_to_fpga:avalonmm_write_slave_write
	wire   [31:0] mm_interconnect_1_fifo_hps_to_fpga_in_writedata;                      // mm_interconnect_1:fifo_hps_to_fpga_in_writedata -> fifo_hps_to_fpga:avalonmm_write_slave_writedata
	wire   [31:0] mm_interconnect_1_fifo_fpga_to_hps_out_readdata;                      // fifo_fpga_to_hps:avalonmm_read_slave_readdata -> mm_interconnect_1:fifo_fpga_to_hps_out_readdata
	wire          mm_interconnect_1_fifo_fpga_to_hps_out_waitrequest;                   // fifo_fpga_to_hps:avalonmm_read_slave_waitrequest -> mm_interconnect_1:fifo_fpga_to_hps_out_waitrequest
	wire          mm_interconnect_1_fifo_fpga_to_hps_out_read;                          // mm_interconnect_1:fifo_fpga_to_hps_out_read -> fifo_fpga_to_hps:avalonmm_read_slave_read
	wire          mm_interconnect_1_ram_s1_chipselect;                                  // mm_interconnect_1:ram_s1_chipselect -> ram:chipselect
	wire   [31:0] mm_interconnect_1_ram_s1_readdata;                                    // ram:readdata -> mm_interconnect_1:ram_s1_readdata
	wire   [10:0] mm_interconnect_1_ram_s1_address;                                     // mm_interconnect_1:ram_s1_address -> ram:address
	wire    [3:0] mm_interconnect_1_ram_s1_byteenable;                                  // mm_interconnect_1:ram_s1_byteenable -> ram:byteenable
	wire          mm_interconnect_1_ram_s1_write;                                       // mm_interconnect_1:ram_s1_write -> ram:write
	wire   [31:0] mm_interconnect_1_ram_s1_writedata;                                   // mm_interconnect_1:ram_s1_writedata -> ram:writedata
	wire          mm_interconnect_1_ram_s1_clken;                                       // mm_interconnect_1:ram_s1_clken -> ram:clken
	wire          mm_interconnect_1_new_sdram_controller_0_s1_chipselect;               // mm_interconnect_1:new_sdram_controller_0_s1_chipselect -> new_sdram_controller_0:az_cs
	wire   [15:0] mm_interconnect_1_new_sdram_controller_0_s1_readdata;                 // new_sdram_controller_0:za_data -> mm_interconnect_1:new_sdram_controller_0_s1_readdata
	wire          mm_interconnect_1_new_sdram_controller_0_s1_waitrequest;              // new_sdram_controller_0:za_waitrequest -> mm_interconnect_1:new_sdram_controller_0_s1_waitrequest
	wire   [24:0] mm_interconnect_1_new_sdram_controller_0_s1_address;                  // mm_interconnect_1:new_sdram_controller_0_s1_address -> new_sdram_controller_0:az_addr
	wire          mm_interconnect_1_new_sdram_controller_0_s1_read;                     // mm_interconnect_1:new_sdram_controller_0_s1_read -> new_sdram_controller_0:az_rd_n
	wire    [1:0] mm_interconnect_1_new_sdram_controller_0_s1_byteenable;               // mm_interconnect_1:new_sdram_controller_0_s1_byteenable -> new_sdram_controller_0:az_be_n
	wire          mm_interconnect_1_new_sdram_controller_0_s1_readdatavalid;            // new_sdram_controller_0:za_valid -> mm_interconnect_1:new_sdram_controller_0_s1_readdatavalid
	wire          mm_interconnect_1_new_sdram_controller_0_s1_write;                    // mm_interconnect_1:new_sdram_controller_0_s1_write -> new_sdram_controller_0:az_wr_n
	wire   [15:0] mm_interconnect_1_new_sdram_controller_0_s1_writedata;                // mm_interconnect_1:new_sdram_controller_0_s1_writedata -> new_sdram_controller_0:az_data
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_awburst;                                 // Arm_A9_HPS:h2f_lw_AWBURST -> mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_awburst
	wire    [3:0] arm_a9_hps_h2f_lw_axi_master_arlen;                                   // Arm_A9_HPS:h2f_lw_ARLEN -> mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_arlen
	wire    [3:0] arm_a9_hps_h2f_lw_axi_master_wstrb;                                   // Arm_A9_HPS:h2f_lw_WSTRB -> mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_wstrb
	wire          arm_a9_hps_h2f_lw_axi_master_wready;                                  // mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_wready -> Arm_A9_HPS:h2f_lw_WREADY
	wire   [11:0] arm_a9_hps_h2f_lw_axi_master_rid;                                     // mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_rid -> Arm_A9_HPS:h2f_lw_RID
	wire          arm_a9_hps_h2f_lw_axi_master_rready;                                  // Arm_A9_HPS:h2f_lw_RREADY -> mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_rready
	wire    [3:0] arm_a9_hps_h2f_lw_axi_master_awlen;                                   // Arm_A9_HPS:h2f_lw_AWLEN -> mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_awlen
	wire   [11:0] arm_a9_hps_h2f_lw_axi_master_wid;                                     // Arm_A9_HPS:h2f_lw_WID -> mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_wid
	wire    [3:0] arm_a9_hps_h2f_lw_axi_master_arcache;                                 // Arm_A9_HPS:h2f_lw_ARCACHE -> mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_arcache
	wire          arm_a9_hps_h2f_lw_axi_master_wvalid;                                  // Arm_A9_HPS:h2f_lw_WVALID -> mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_wvalid
	wire   [20:0] arm_a9_hps_h2f_lw_axi_master_araddr;                                  // Arm_A9_HPS:h2f_lw_ARADDR -> mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_araddr
	wire    [2:0] arm_a9_hps_h2f_lw_axi_master_arprot;                                  // Arm_A9_HPS:h2f_lw_ARPROT -> mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_arprot
	wire    [2:0] arm_a9_hps_h2f_lw_axi_master_awprot;                                  // Arm_A9_HPS:h2f_lw_AWPROT -> mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_awprot
	wire   [31:0] arm_a9_hps_h2f_lw_axi_master_wdata;                                   // Arm_A9_HPS:h2f_lw_WDATA -> mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_wdata
	wire          arm_a9_hps_h2f_lw_axi_master_arvalid;                                 // Arm_A9_HPS:h2f_lw_ARVALID -> mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_arvalid
	wire    [3:0] arm_a9_hps_h2f_lw_axi_master_awcache;                                 // Arm_A9_HPS:h2f_lw_AWCACHE -> mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_awcache
	wire   [11:0] arm_a9_hps_h2f_lw_axi_master_arid;                                    // Arm_A9_HPS:h2f_lw_ARID -> mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_arid
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_arlock;                                  // Arm_A9_HPS:h2f_lw_ARLOCK -> mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_arlock
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_awlock;                                  // Arm_A9_HPS:h2f_lw_AWLOCK -> mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_awlock
	wire   [20:0] arm_a9_hps_h2f_lw_axi_master_awaddr;                                  // Arm_A9_HPS:h2f_lw_AWADDR -> mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_awaddr
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_bresp;                                   // mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_bresp -> Arm_A9_HPS:h2f_lw_BRESP
	wire          arm_a9_hps_h2f_lw_axi_master_arready;                                 // mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_arready -> Arm_A9_HPS:h2f_lw_ARREADY
	wire   [31:0] arm_a9_hps_h2f_lw_axi_master_rdata;                                   // mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_rdata -> Arm_A9_HPS:h2f_lw_RDATA
	wire          arm_a9_hps_h2f_lw_axi_master_awready;                                 // mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_awready -> Arm_A9_HPS:h2f_lw_AWREADY
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_arburst;                                 // Arm_A9_HPS:h2f_lw_ARBURST -> mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_arburst
	wire    [2:0] arm_a9_hps_h2f_lw_axi_master_arsize;                                  // Arm_A9_HPS:h2f_lw_ARSIZE -> mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_arsize
	wire          arm_a9_hps_h2f_lw_axi_master_bready;                                  // Arm_A9_HPS:h2f_lw_BREADY -> mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_bready
	wire          arm_a9_hps_h2f_lw_axi_master_rlast;                                   // mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_rlast -> Arm_A9_HPS:h2f_lw_RLAST
	wire          arm_a9_hps_h2f_lw_axi_master_wlast;                                   // Arm_A9_HPS:h2f_lw_WLAST -> mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_wlast
	wire    [1:0] arm_a9_hps_h2f_lw_axi_master_rresp;                                   // mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_rresp -> Arm_A9_HPS:h2f_lw_RRESP
	wire   [11:0] arm_a9_hps_h2f_lw_axi_master_awid;                                    // Arm_A9_HPS:h2f_lw_AWID -> mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_awid
	wire   [11:0] arm_a9_hps_h2f_lw_axi_master_bid;                                     // mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_bid -> Arm_A9_HPS:h2f_lw_BID
	wire          arm_a9_hps_h2f_lw_axi_master_bvalid;                                  // mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_bvalid -> Arm_A9_HPS:h2f_lw_BVALID
	wire    [2:0] arm_a9_hps_h2f_lw_axi_master_awsize;                                  // Arm_A9_HPS:h2f_lw_AWSIZE -> mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_awsize
	wire          arm_a9_hps_h2f_lw_axi_master_awvalid;                                 // Arm_A9_HPS:h2f_lw_AWVALID -> mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_awvalid
	wire          arm_a9_hps_h2f_lw_axi_master_rvalid;                                  // mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_rvalid -> Arm_A9_HPS:h2f_lw_RVALID
	wire          mm_interconnect_2_system_console_avalon_jtag_slave_chipselect;        // mm_interconnect_2:system_console_avalon_jtag_slave_chipselect -> system_console:av_chipselect
	wire   [31:0] mm_interconnect_2_system_console_avalon_jtag_slave_readdata;          // system_console:av_readdata -> mm_interconnect_2:system_console_avalon_jtag_slave_readdata
	wire          mm_interconnect_2_system_console_avalon_jtag_slave_waitrequest;       // system_console:av_waitrequest -> mm_interconnect_2:system_console_avalon_jtag_slave_waitrequest
	wire    [0:0] mm_interconnect_2_system_console_avalon_jtag_slave_address;           // mm_interconnect_2:system_console_avalon_jtag_slave_address -> system_console:av_address
	wire          mm_interconnect_2_system_console_avalon_jtag_slave_read;              // mm_interconnect_2:system_console_avalon_jtag_slave_read -> system_console:av_read_n
	wire          mm_interconnect_2_system_console_avalon_jtag_slave_write;             // mm_interconnect_2:system_console_avalon_jtag_slave_write -> system_console:av_write_n
	wire   [31:0] mm_interconnect_2_system_console_avalon_jtag_slave_writedata;         // mm_interconnect_2:system_console_avalon_jtag_slave_writedata -> system_console:av_writedata
	wire   [31:0] mm_interconnect_2_alt_vip_vfr_0_avalon_slave_readdata;                // alt_vip_vfr_0:slave_readdata -> mm_interconnect_2:alt_vip_vfr_0_avalon_slave_readdata
	wire    [4:0] mm_interconnect_2_alt_vip_vfr_0_avalon_slave_address;                 // mm_interconnect_2:alt_vip_vfr_0_avalon_slave_address -> alt_vip_vfr_0:slave_address
	wire          mm_interconnect_2_alt_vip_vfr_0_avalon_slave_read;                    // mm_interconnect_2:alt_vip_vfr_0_avalon_slave_read -> alt_vip_vfr_0:slave_read
	wire          mm_interconnect_2_alt_vip_vfr_0_avalon_slave_write;                   // mm_interconnect_2:alt_vip_vfr_0_avalon_slave_write -> alt_vip_vfr_0:slave_write
	wire   [31:0] mm_interconnect_2_alt_vip_vfr_0_avalon_slave_writedata;               // mm_interconnect_2:alt_vip_vfr_0_avalon_slave_writedata -> alt_vip_vfr_0:slave_writedata
	wire          mm_interconnect_2_reg32_avalon_interface_0_avalon_slave_0_chipselect; // mm_interconnect_2:reg32_avalon_interface_0_avalon_slave_0_chipselect -> reg32_avalon_interface_0:chipselect
	wire   [31:0] mm_interconnect_2_reg32_avalon_interface_0_avalon_slave_0_readdata;   // reg32_avalon_interface_0:readdata -> mm_interconnect_2:reg32_avalon_interface_0_avalon_slave_0_readdata
	wire          mm_interconnect_2_reg32_avalon_interface_0_avalon_slave_0_read;       // mm_interconnect_2:reg32_avalon_interface_0_avalon_slave_0_read -> reg32_avalon_interface_0:read
	wire    [3:0] mm_interconnect_2_reg32_avalon_interface_0_avalon_slave_0_byteenable; // mm_interconnect_2:reg32_avalon_interface_0_avalon_slave_0_byteenable -> reg32_avalon_interface_0:byteenable
	wire          mm_interconnect_2_reg32_avalon_interface_0_avalon_slave_0_write;      // mm_interconnect_2:reg32_avalon_interface_0_avalon_slave_0_write -> reg32_avalon_interface_0:write
	wire   [31:0] mm_interconnect_2_reg32_avalon_interface_0_avalon_slave_0_writedata;  // mm_interconnect_2:reg32_avalon_interface_0_avalon_slave_0_writedata -> reg32_avalon_interface_0:writedata
	wire   [31:0] mm_interconnect_2_sysid_qsys_0_control_slave_readdata;                // sysid_qsys_0:readdata -> mm_interconnect_2:sysid_qsys_0_control_slave_readdata
	wire    [0:0] mm_interconnect_2_sysid_qsys_0_control_slave_address;                 // mm_interconnect_2:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire   [31:0] mm_interconnect_2_fifo_hps_to_fpga_in_csr_readdata;                   // fifo_hps_to_fpga:wrclk_control_slave_readdata -> mm_interconnect_2:fifo_hps_to_fpga_in_csr_readdata
	wire    [2:0] mm_interconnect_2_fifo_hps_to_fpga_in_csr_address;                    // mm_interconnect_2:fifo_hps_to_fpga_in_csr_address -> fifo_hps_to_fpga:wrclk_control_slave_address
	wire          mm_interconnect_2_fifo_hps_to_fpga_in_csr_read;                       // mm_interconnect_2:fifo_hps_to_fpga_in_csr_read -> fifo_hps_to_fpga:wrclk_control_slave_read
	wire          mm_interconnect_2_fifo_hps_to_fpga_in_csr_write;                      // mm_interconnect_2:fifo_hps_to_fpga_in_csr_write -> fifo_hps_to_fpga:wrclk_control_slave_write
	wire   [31:0] mm_interconnect_2_fifo_hps_to_fpga_in_csr_writedata;                  // mm_interconnect_2:fifo_hps_to_fpga_in_csr_writedata -> fifo_hps_to_fpga:wrclk_control_slave_writedata
	wire   [31:0] mm_interconnect_2_fifo_fpga_to_hps_out_csr_readdata;                  // fifo_fpga_to_hps:rdclk_control_slave_readdata -> mm_interconnect_2:fifo_fpga_to_hps_out_csr_readdata
	wire    [2:0] mm_interconnect_2_fifo_fpga_to_hps_out_csr_address;                   // mm_interconnect_2:fifo_fpga_to_hps_out_csr_address -> fifo_fpga_to_hps:rdclk_control_slave_address
	wire          mm_interconnect_2_fifo_fpga_to_hps_out_csr_read;                      // mm_interconnect_2:fifo_fpga_to_hps_out_csr_read -> fifo_fpga_to_hps:rdclk_control_slave_read
	wire          mm_interconnect_2_fifo_fpga_to_hps_out_csr_write;                     // mm_interconnect_2:fifo_fpga_to_hps_out_csr_write -> fifo_fpga_to_hps:rdclk_control_slave_write
	wire   [31:0] mm_interconnect_2_fifo_fpga_to_hps_out_csr_writedata;                 // mm_interconnect_2:fifo_fpga_to_hps_out_csr_writedata -> fifo_fpga_to_hps:rdclk_control_slave_writedata
	wire          mm_interconnect_2_hex5_hex0_s1_chipselect;                            // mm_interconnect_2:hex5_hex0_s1_chipselect -> hex5_hex0:chipselect
	wire   [31:0] mm_interconnect_2_hex5_hex0_s1_readdata;                              // hex5_hex0:readdata -> mm_interconnect_2:hex5_hex0_s1_readdata
	wire    [1:0] mm_interconnect_2_hex5_hex0_s1_address;                               // mm_interconnect_2:hex5_hex0_s1_address -> hex5_hex0:address
	wire          mm_interconnect_2_hex5_hex0_s1_write;                                 // mm_interconnect_2:hex5_hex0_s1_write -> hex5_hex0:write_n
	wire   [31:0] mm_interconnect_2_hex5_hex0_s1_writedata;                             // mm_interconnect_2:hex5_hex0_s1_writedata -> hex5_hex0:writedata
	wire          mm_interconnect_2_pushbuttons_s1_chipselect;                          // mm_interconnect_2:pushbuttons_s1_chipselect -> pushbuttons:chipselect
	wire   [31:0] mm_interconnect_2_pushbuttons_s1_readdata;                            // pushbuttons:readdata -> mm_interconnect_2:pushbuttons_s1_readdata
	wire    [1:0] mm_interconnect_2_pushbuttons_s1_address;                             // mm_interconnect_2:pushbuttons_s1_address -> pushbuttons:address
	wire          mm_interconnect_2_pushbuttons_s1_write;                               // mm_interconnect_2:pushbuttons_s1_write -> pushbuttons:write_n
	wire   [31:0] mm_interconnect_2_pushbuttons_s1_writedata;                           // mm_interconnect_2:pushbuttons_s1_writedata -> pushbuttons:writedata
	wire          irq_mapper_receiver0_irq;                                             // system_console:av_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                             // pushbuttons:irq -> irq_mapper:receiver1_irq
	wire   [31:0] arm_a9_hps_f2h_irq0_irq;                                              // irq_mapper:sender_irq -> Arm_A9_HPS:f2h_irq_p0
	wire   [31:0] arm_a9_hps_f2h_irq1_irq;                                              // irq_mapper_001:sender_irq -> Arm_A9_HPS:f2h_irq_p1
	wire          rst_controller_reset_out_reset;                                       // rst_controller:reset_out -> [alt_vip_itc_0:rst, alt_vip_vfr_0:reset, mm_interconnect_2:alt_vip_vfr_0_clock_reset_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_001_reset_out_reset;                                   // rst_controller_001:reset_out -> [alt_vip_vfr_0:master_reset, mm_interconnect_0:alt_vip_vfr_0_clock_master_reset_reset_bridge_in_reset_reset, mm_interconnect_2:sysid_qsys_0_reset_reset_bridge_in_reset_reset, sysid_qsys_0:reset_n]
	wire          rst_controller_002_reset_out_reset;                                   // rst_controller_002:reset_out -> [fifo_fpga_to_hps:wrreset_n, fifo_hps_to_fpga:rdreset_n, ram:reset2]
	wire          rst_controller_002_reset_out_reset_req;                               // rst_controller_002:reset_req -> [ram:reset_req2, rst_translator:reset_req_in]
	wire          arm_a9_hps_h2f_reset_reset;                                           // Arm_A9_HPS:h2f_rst_n -> [rst_controller_002:reset_in0, rst_controller_003:reset_in0, rst_controller_004:reset_in0]
	wire          rst_controller_003_reset_out_reset;                                   // rst_controller_003:reset_out -> [fifo_fpga_to_hps:rdreset_n, fifo_hps_to_fpga:wrreset_n, hex5_hex0:reset_n, mm_interconnect_1:fifo_hps_to_fpga_reset_in_reset_bridge_in_reset_reset, mm_interconnect_2:system_console_reset_reset_bridge_in_reset_reset, new_sdram_controller_0:reset_n, pushbuttons:reset_n, ram:reset, reg32_avalon_interface_0:reset_n, rst_translator_001:in_reset, system_console:rst_n]
	wire          rst_controller_003_reset_out_reset_req;                               // rst_controller_003:reset_req -> [ram:reset_req, rst_translator_001:reset_req_in]
	wire          rst_controller_004_reset_out_reset;                                   // rst_controller_004:reset_out -> [mm_interconnect_0:Arm_A9_HPS_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:Arm_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_2:Arm_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]

	sys_vga_Arm_A9_HPS #(
		.F2S_Width (2),
		.S2F_Width (3)
	) arm_a9_hps (
		.f2h_boot_from_fpga_ready      (),                                                   // f2h_boot_from_fpga.boot_from_fpga_ready
		.f2h_boot_from_fpga_on_failure (),                                                   //                   .boot_from_fpga_on_failure
		.mem_a                         (memory_mem_a),                                       //             memory.mem_a
		.mem_ba                        (memory_mem_ba),                                      //                   .mem_ba
		.mem_ck                        (memory_mem_ck),                                      //                   .mem_ck
		.mem_ck_n                      (memory_mem_ck_n),                                    //                   .mem_ck_n
		.mem_cke                       (memory_mem_cke),                                     //                   .mem_cke
		.mem_cs_n                      (memory_mem_cs_n),                                    //                   .mem_cs_n
		.mem_ras_n                     (memory_mem_ras_n),                                   //                   .mem_ras_n
		.mem_cas_n                     (memory_mem_cas_n),                                   //                   .mem_cas_n
		.mem_we_n                      (memory_mem_we_n),                                    //                   .mem_we_n
		.mem_reset_n                   (memory_mem_reset_n),                                 //                   .mem_reset_n
		.mem_dq                        (memory_mem_dq),                                      //                   .mem_dq
		.mem_dqs                       (memory_mem_dqs),                                     //                   .mem_dqs
		.mem_dqs_n                     (memory_mem_dqs_n),                                   //                   .mem_dqs_n
		.mem_odt                       (memory_mem_odt),                                     //                   .mem_odt
		.mem_dm                        (memory_mem_dm),                                      //                   .mem_dm
		.oct_rzqin                     (memory_oct_rzqin),                                   //                   .oct_rzqin
		.hps_io_sdio_inst_CMD          (hps_io_hps_io_sdio_inst_CMD),                        //             hps_io.hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0           (hps_io_hps_io_sdio_inst_D0),                         //                   .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1           (hps_io_hps_io_sdio_inst_D1),                         //                   .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK          (hps_io_hps_io_sdio_inst_CLK),                        //                   .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2           (hps_io_hps_io_sdio_inst_D2),                         //                   .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3           (hps_io_hps_io_sdio_inst_D3),                         //                   .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0           (hps_io_hps_io_usb1_inst_D0),                         //                   .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1           (hps_io_hps_io_usb1_inst_D1),                         //                   .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2           (hps_io_hps_io_usb1_inst_D2),                         //                   .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3           (hps_io_hps_io_usb1_inst_D3),                         //                   .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4           (hps_io_hps_io_usb1_inst_D4),                         //                   .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5           (hps_io_hps_io_usb1_inst_D5),                         //                   .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6           (hps_io_hps_io_usb1_inst_D6),                         //                   .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7           (hps_io_hps_io_usb1_inst_D7),                         //                   .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK          (hps_io_hps_io_usb1_inst_CLK),                        //                   .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP          (hps_io_hps_io_usb1_inst_STP),                        //                   .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR          (hps_io_hps_io_usb1_inst_DIR),                        //                   .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT          (hps_io_hps_io_usb1_inst_NXT),                        //                   .hps_io_usb1_inst_NXT
		.hps_io_uart0_inst_RX          (hps_io_hps_io_uart0_inst_RX),                        //                   .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX          (hps_io_hps_io_uart0_inst_TX),                        //                   .hps_io_uart0_inst_TX
		.h2f_rst_n                     (arm_a9_hps_h2f_reset_reset),                         //          h2f_reset.reset_n
		.h2f_axi_clk                   (sys_sdram_pll_0_sys_clk_clk),                        //      h2f_axi_clock.clk
		.h2f_AWID                      (arm_a9_hps_h2f_axi_master_awid),                     //     h2f_axi_master.awid
		.h2f_AWADDR                    (arm_a9_hps_h2f_axi_master_awaddr),                   //                   .awaddr
		.h2f_AWLEN                     (arm_a9_hps_h2f_axi_master_awlen),                    //                   .awlen
		.h2f_AWSIZE                    (arm_a9_hps_h2f_axi_master_awsize),                   //                   .awsize
		.h2f_AWBURST                   (arm_a9_hps_h2f_axi_master_awburst),                  //                   .awburst
		.h2f_AWLOCK                    (arm_a9_hps_h2f_axi_master_awlock),                   //                   .awlock
		.h2f_AWCACHE                   (arm_a9_hps_h2f_axi_master_awcache),                  //                   .awcache
		.h2f_AWPROT                    (arm_a9_hps_h2f_axi_master_awprot),                   //                   .awprot
		.h2f_AWVALID                   (arm_a9_hps_h2f_axi_master_awvalid),                  //                   .awvalid
		.h2f_AWREADY                   (arm_a9_hps_h2f_axi_master_awready),                  //                   .awready
		.h2f_WID                       (arm_a9_hps_h2f_axi_master_wid),                      //                   .wid
		.h2f_WDATA                     (arm_a9_hps_h2f_axi_master_wdata),                    //                   .wdata
		.h2f_WSTRB                     (arm_a9_hps_h2f_axi_master_wstrb),                    //                   .wstrb
		.h2f_WLAST                     (arm_a9_hps_h2f_axi_master_wlast),                    //                   .wlast
		.h2f_WVALID                    (arm_a9_hps_h2f_axi_master_wvalid),                   //                   .wvalid
		.h2f_WREADY                    (arm_a9_hps_h2f_axi_master_wready),                   //                   .wready
		.h2f_BID                       (arm_a9_hps_h2f_axi_master_bid),                      //                   .bid
		.h2f_BRESP                     (arm_a9_hps_h2f_axi_master_bresp),                    //                   .bresp
		.h2f_BVALID                    (arm_a9_hps_h2f_axi_master_bvalid),                   //                   .bvalid
		.h2f_BREADY                    (arm_a9_hps_h2f_axi_master_bready),                   //                   .bready
		.h2f_ARID                      (arm_a9_hps_h2f_axi_master_arid),                     //                   .arid
		.h2f_ARADDR                    (arm_a9_hps_h2f_axi_master_araddr),                   //                   .araddr
		.h2f_ARLEN                     (arm_a9_hps_h2f_axi_master_arlen),                    //                   .arlen
		.h2f_ARSIZE                    (arm_a9_hps_h2f_axi_master_arsize),                   //                   .arsize
		.h2f_ARBURST                   (arm_a9_hps_h2f_axi_master_arburst),                  //                   .arburst
		.h2f_ARLOCK                    (arm_a9_hps_h2f_axi_master_arlock),                   //                   .arlock
		.h2f_ARCACHE                   (arm_a9_hps_h2f_axi_master_arcache),                  //                   .arcache
		.h2f_ARPROT                    (arm_a9_hps_h2f_axi_master_arprot),                   //                   .arprot
		.h2f_ARVALID                   (arm_a9_hps_h2f_axi_master_arvalid),                  //                   .arvalid
		.h2f_ARREADY                   (arm_a9_hps_h2f_axi_master_arready),                  //                   .arready
		.h2f_RID                       (arm_a9_hps_h2f_axi_master_rid),                      //                   .rid
		.h2f_RDATA                     (arm_a9_hps_h2f_axi_master_rdata),                    //                   .rdata
		.h2f_RRESP                     (arm_a9_hps_h2f_axi_master_rresp),                    //                   .rresp
		.h2f_RLAST                     (arm_a9_hps_h2f_axi_master_rlast),                    //                   .rlast
		.h2f_RVALID                    (arm_a9_hps_h2f_axi_master_rvalid),                   //                   .rvalid
		.h2f_RREADY                    (arm_a9_hps_h2f_axi_master_rready),                   //                   .rready
		.f2h_axi_clk                   (sys_sdram_pll_0_sys_clk_clk),                        //      f2h_axi_clock.clk
		.f2h_AWID                      (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awid),    //      f2h_axi_slave.awid
		.f2h_AWADDR                    (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awaddr),  //                   .awaddr
		.f2h_AWLEN                     (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awlen),   //                   .awlen
		.f2h_AWSIZE                    (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awsize),  //                   .awsize
		.f2h_AWBURST                   (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awburst), //                   .awburst
		.f2h_AWLOCK                    (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awlock),  //                   .awlock
		.f2h_AWCACHE                   (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awcache), //                   .awcache
		.f2h_AWPROT                    (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awprot),  //                   .awprot
		.f2h_AWVALID                   (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awvalid), //                   .awvalid
		.f2h_AWREADY                   (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awready), //                   .awready
		.f2h_AWUSER                    (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awuser),  //                   .awuser
		.f2h_WID                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wid),     //                   .wid
		.f2h_WDATA                     (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wdata),   //                   .wdata
		.f2h_WSTRB                     (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wstrb),   //                   .wstrb
		.f2h_WLAST                     (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wlast),   //                   .wlast
		.f2h_WVALID                    (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wvalid),  //                   .wvalid
		.f2h_WREADY                    (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wready),  //                   .wready
		.f2h_BID                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bid),     //                   .bid
		.f2h_BRESP                     (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bresp),   //                   .bresp
		.f2h_BVALID                    (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bvalid),  //                   .bvalid
		.f2h_BREADY                    (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bready),  //                   .bready
		.f2h_ARID                      (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arid),    //                   .arid
		.f2h_ARADDR                    (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_araddr),  //                   .araddr
		.f2h_ARLEN                     (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arlen),   //                   .arlen
		.f2h_ARSIZE                    (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arsize),  //                   .arsize
		.f2h_ARBURST                   (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arburst), //                   .arburst
		.f2h_ARLOCK                    (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arlock),  //                   .arlock
		.f2h_ARCACHE                   (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arcache), //                   .arcache
		.f2h_ARPROT                    (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arprot),  //                   .arprot
		.f2h_ARVALID                   (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arvalid), //                   .arvalid
		.f2h_ARREADY                   (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arready), //                   .arready
		.f2h_ARUSER                    (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_aruser),  //                   .aruser
		.f2h_RID                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rid),     //                   .rid
		.f2h_RDATA                     (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rdata),   //                   .rdata
		.f2h_RRESP                     (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rresp),   //                   .rresp
		.f2h_RLAST                     (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rlast),   //                   .rlast
		.f2h_RVALID                    (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rvalid),  //                   .rvalid
		.f2h_RREADY                    (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rready),  //                   .rready
		.h2f_lw_axi_clk                (sys_sdram_pll_0_sys_clk_clk),                        //   h2f_lw_axi_clock.clk
		.h2f_lw_AWID                   (arm_a9_hps_h2f_lw_axi_master_awid),                  //  h2f_lw_axi_master.awid
		.h2f_lw_AWADDR                 (arm_a9_hps_h2f_lw_axi_master_awaddr),                //                   .awaddr
		.h2f_lw_AWLEN                  (arm_a9_hps_h2f_lw_axi_master_awlen),                 //                   .awlen
		.h2f_lw_AWSIZE                 (arm_a9_hps_h2f_lw_axi_master_awsize),                //                   .awsize
		.h2f_lw_AWBURST                (arm_a9_hps_h2f_lw_axi_master_awburst),               //                   .awburst
		.h2f_lw_AWLOCK                 (arm_a9_hps_h2f_lw_axi_master_awlock),                //                   .awlock
		.h2f_lw_AWCACHE                (arm_a9_hps_h2f_lw_axi_master_awcache),               //                   .awcache
		.h2f_lw_AWPROT                 (arm_a9_hps_h2f_lw_axi_master_awprot),                //                   .awprot
		.h2f_lw_AWVALID                (arm_a9_hps_h2f_lw_axi_master_awvalid),               //                   .awvalid
		.h2f_lw_AWREADY                (arm_a9_hps_h2f_lw_axi_master_awready),               //                   .awready
		.h2f_lw_WID                    (arm_a9_hps_h2f_lw_axi_master_wid),                   //                   .wid
		.h2f_lw_WDATA                  (arm_a9_hps_h2f_lw_axi_master_wdata),                 //                   .wdata
		.h2f_lw_WSTRB                  (arm_a9_hps_h2f_lw_axi_master_wstrb),                 //                   .wstrb
		.h2f_lw_WLAST                  (arm_a9_hps_h2f_lw_axi_master_wlast),                 //                   .wlast
		.h2f_lw_WVALID                 (arm_a9_hps_h2f_lw_axi_master_wvalid),                //                   .wvalid
		.h2f_lw_WREADY                 (arm_a9_hps_h2f_lw_axi_master_wready),                //                   .wready
		.h2f_lw_BID                    (arm_a9_hps_h2f_lw_axi_master_bid),                   //                   .bid
		.h2f_lw_BRESP                  (arm_a9_hps_h2f_lw_axi_master_bresp),                 //                   .bresp
		.h2f_lw_BVALID                 (arm_a9_hps_h2f_lw_axi_master_bvalid),                //                   .bvalid
		.h2f_lw_BREADY                 (arm_a9_hps_h2f_lw_axi_master_bready),                //                   .bready
		.h2f_lw_ARID                   (arm_a9_hps_h2f_lw_axi_master_arid),                  //                   .arid
		.h2f_lw_ARADDR                 (arm_a9_hps_h2f_lw_axi_master_araddr),                //                   .araddr
		.h2f_lw_ARLEN                  (arm_a9_hps_h2f_lw_axi_master_arlen),                 //                   .arlen
		.h2f_lw_ARSIZE                 (arm_a9_hps_h2f_lw_axi_master_arsize),                //                   .arsize
		.h2f_lw_ARBURST                (arm_a9_hps_h2f_lw_axi_master_arburst),               //                   .arburst
		.h2f_lw_ARLOCK                 (arm_a9_hps_h2f_lw_axi_master_arlock),                //                   .arlock
		.h2f_lw_ARCACHE                (arm_a9_hps_h2f_lw_axi_master_arcache),               //                   .arcache
		.h2f_lw_ARPROT                 (arm_a9_hps_h2f_lw_axi_master_arprot),                //                   .arprot
		.h2f_lw_ARVALID                (arm_a9_hps_h2f_lw_axi_master_arvalid),               //                   .arvalid
		.h2f_lw_ARREADY                (arm_a9_hps_h2f_lw_axi_master_arready),               //                   .arready
		.h2f_lw_RID                    (arm_a9_hps_h2f_lw_axi_master_rid),                   //                   .rid
		.h2f_lw_RDATA                  (arm_a9_hps_h2f_lw_axi_master_rdata),                 //                   .rdata
		.h2f_lw_RRESP                  (arm_a9_hps_h2f_lw_axi_master_rresp),                 //                   .rresp
		.h2f_lw_RLAST                  (arm_a9_hps_h2f_lw_axi_master_rlast),                 //                   .rlast
		.h2f_lw_RVALID                 (arm_a9_hps_h2f_lw_axi_master_rvalid),                //                   .rvalid
		.h2f_lw_RREADY                 (arm_a9_hps_h2f_lw_axi_master_rready),                //                   .rready
		.f2h_irq_p0                    (arm_a9_hps_f2h_irq0_irq),                            //           f2h_irq0.irq
		.f2h_irq_p1                    (arm_a9_hps_f2h_irq1_irq)                             //           f2h_irq1.irq
	);

	alt_vipitc131_IS2Vid #(
		.NUMBER_OF_COLOUR_PLANES       (4),
		.COLOUR_PLANES_ARE_IN_PARALLEL (1),
		.BPS                           (8),
		.INTERLACED                    (0),
		.H_ACTIVE_PIXELS               (1024),
		.V_ACTIVE_LINES                (768),
		.ACCEPT_COLOURS_IN_SEQ         (0),
		.FIFO_DEPTH                    (1920),
		.CLOCKS_ARE_SAME               (0),
		.USE_CONTROL                   (0),
		.NO_OF_MODES                   (1),
		.THRESHOLD                     (1919),
		.STD_WIDTH                     (1),
		.GENERATE_SYNC                 (0),
		.USE_EMBEDDED_SYNCS            (0),
		.AP_LINE                       (0),
		.V_BLANK                       (0),
		.H_BLANK                       (0),
		.H_SYNC_LENGTH                 (136),
		.H_FRONT_PORCH                 (24),
		.H_BACK_PORCH                  (160),
		.V_SYNC_LENGTH                 (6),
		.V_FRONT_PORCH                 (3),
		.V_BACK_PORCH                  (29),
		.F_RISING_EDGE                 (0),
		.F_FALLING_EDGE                (0),
		.FIELD0_V_RISING_EDGE          (0),
		.FIELD0_V_BLANK                (0),
		.FIELD0_V_SYNC_LENGTH          (0),
		.FIELD0_V_FRONT_PORCH          (0),
		.FIELD0_V_BACK_PORCH           (0),
		.ANC_LINE                      (0),
		.FIELD0_ANC_LINE               (0)
	) alt_vip_itc_0 (
		.is_clk        (pll_0_outclk0_clk),                                   //       is_clk_rst.clk
		.rst           (rst_controller_reset_out_reset),                      // is_clk_rst_reset.reset
		.is_data       (alt_vip_vfr_0_avalon_streaming_source_data),          //              din.data
		.is_valid      (alt_vip_vfr_0_avalon_streaming_source_valid),         //                 .valid
		.is_ready      (alt_vip_vfr_0_avalon_streaming_source_ready),         //                 .ready
		.is_sop        (alt_vip_vfr_0_avalon_streaming_source_startofpacket), //                 .startofpacket
		.is_eop        (alt_vip_vfr_0_avalon_streaming_source_endofpacket),   //                 .endofpacket
		.vid_clk       (alt_vip_itc_0_clocked_video_vid_clk),                 //    clocked_video.export
		.vid_data      (alt_vip_itc_0_clocked_video_vid_data),                //                 .export
		.underflow     (alt_vip_itc_0_clocked_video_underflow),               //                 .export
		.vid_datavalid (alt_vip_itc_0_clocked_video_vid_datavalid),           //                 .export
		.vid_v_sync    (alt_vip_itc_0_clocked_video_vid_v_sync),              //                 .export
		.vid_h_sync    (alt_vip_itc_0_clocked_video_vid_h_sync),              //                 .export
		.vid_f         (alt_vip_itc_0_clocked_video_vid_f),                   //                 .export
		.vid_h         (alt_vip_itc_0_clocked_video_vid_h),                   //                 .export
		.vid_v         (alt_vip_itc_0_clocked_video_vid_v)                    //                 .export
	);

	sys_vga_alt_vip_vfr_0 alt_vip_vfr_0 (
		.clock                (pll_0_outclk0_clk),                                      //             clock_reset.clk
		.reset                (rst_controller_reset_out_reset),                         //       clock_reset_reset.reset
		.master_clock         (sys_sdram_pll_0_sys_clk_clk),                            //            clock_master.clk
		.master_reset         (rst_controller_001_reset_out_reset),                     //      clock_master_reset.reset
		.slave_address        (mm_interconnect_2_alt_vip_vfr_0_avalon_slave_address),   //            avalon_slave.address
		.slave_write          (mm_interconnect_2_alt_vip_vfr_0_avalon_slave_write),     //                        .write
		.slave_writedata      (mm_interconnect_2_alt_vip_vfr_0_avalon_slave_writedata), //                        .writedata
		.slave_read           (mm_interconnect_2_alt_vip_vfr_0_avalon_slave_read),      //                        .read
		.slave_readdata       (mm_interconnect_2_alt_vip_vfr_0_avalon_slave_readdata),  //                        .readdata
		.slave_irq            (),                                                       //        interrupt_sender.irq
		.dout_data            (alt_vip_vfr_0_avalon_streaming_source_data),             // avalon_streaming_source.data
		.dout_valid           (alt_vip_vfr_0_avalon_streaming_source_valid),            //                        .valid
		.dout_ready           (alt_vip_vfr_0_avalon_streaming_source_ready),            //                        .ready
		.dout_startofpacket   (alt_vip_vfr_0_avalon_streaming_source_startofpacket),    //                        .startofpacket
		.dout_endofpacket     (alt_vip_vfr_0_avalon_streaming_source_endofpacket),      //                        .endofpacket
		.master_address       (alt_vip_vfr_0_avalon_master_address),                    //           avalon_master.address
		.master_burstcount    (alt_vip_vfr_0_avalon_master_burstcount),                 //                        .burstcount
		.master_readdata      (alt_vip_vfr_0_avalon_master_readdata),                   //                        .readdata
		.master_read          (alt_vip_vfr_0_avalon_master_read),                       //                        .read
		.master_readdatavalid (alt_vip_vfr_0_avalon_master_readdatavalid),              //                        .readdatavalid
		.master_waitrequest   (alt_vip_vfr_0_avalon_master_waitrequest)                 //                        .waitrequest
	);

	sys_vga_fifo_fpga_to_hps fifo_fpga_to_hps (
		.wrclock                          (clock_bridge_0_in_clk_clk),                            //    clk_in.clk
		.wrreset_n                        (~rst_controller_002_reset_out_reset),                  //  reset_in.reset_n
		.rdclock                          (sys_sdram_pll_0_sys_clk_clk),                          //   clk_out.clk
		.rdreset_n                        (~rst_controller_003_reset_out_reset),                  // reset_out.reset_n
		.avalonmm_write_slave_writedata   (fifo_fpga_to_hps_in_writedata),                        //        in.writedata
		.avalonmm_write_slave_write       (fifo_fpga_to_hps_in_write),                            //          .write
		.avalonmm_write_slave_waitrequest (fifo_fpga_to_hps_in_waitrequest),                      //          .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_1_fifo_fpga_to_hps_out_readdata),      //       out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_1_fifo_fpga_to_hps_out_read),          //          .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_1_fifo_fpga_to_hps_out_waitrequest),   //          .waitrequest
		.rdclk_control_slave_address      (mm_interconnect_2_fifo_fpga_to_hps_out_csr_address),   //   out_csr.address
		.rdclk_control_slave_read         (mm_interconnect_2_fifo_fpga_to_hps_out_csr_read),      //          .read
		.rdclk_control_slave_writedata    (mm_interconnect_2_fifo_fpga_to_hps_out_csr_writedata), //          .writedata
		.rdclk_control_slave_write        (mm_interconnect_2_fifo_fpga_to_hps_out_csr_write),     //          .write
		.rdclk_control_slave_readdata     (mm_interconnect_2_fifo_fpga_to_hps_out_csr_readdata),  //          .readdata
		.wrclk_control_slave_address      (fifo_fpga_to_hps_in_csr_address),                      //    in_csr.address
		.wrclk_control_slave_read         (fifo_fpga_to_hps_in_csr_read),                         //          .read
		.wrclk_control_slave_writedata    (fifo_fpga_to_hps_in_csr_writedata),                    //          .writedata
		.wrclk_control_slave_write        (fifo_fpga_to_hps_in_csr_write),                        //          .write
		.wrclk_control_slave_readdata     (fifo_fpga_to_hps_in_csr_readdata)                      //          .readdata
	);

	sys_vga_fifo_fpga_to_hps fifo_hps_to_fpga (
		.wrclock                          (sys_sdram_pll_0_sys_clk_clk),                         //    clk_in.clk
		.wrreset_n                        (~rst_controller_003_reset_out_reset),                 //  reset_in.reset_n
		.rdclock                          (clock_bridge_0_in_clk_clk),                           //   clk_out.clk
		.rdreset_n                        (~rst_controller_002_reset_out_reset),                 // reset_out.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_1_fifo_hps_to_fpga_in_writedata),     //        in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_1_fifo_hps_to_fpga_in_write),         //          .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_1_fifo_hps_to_fpga_in_waitrequest),   //          .waitrequest
		.avalonmm_read_slave_readdata     (fifo_hps_to_fpga_out_readdata),                       //       out.readdata
		.avalonmm_read_slave_read         (fifo_hps_to_fpga_out_read),                           //          .read
		.avalonmm_read_slave_waitrequest  (fifo_hps_to_fpga_out_waitrequest),                    //          .waitrequest
		.rdclk_control_slave_address      (fifo_hps_to_fpga_out_csr_address),                    //   out_csr.address
		.rdclk_control_slave_read         (fifo_hps_to_fpga_out_csr_read),                       //          .read
		.rdclk_control_slave_writedata    (fifo_hps_to_fpga_out_csr_writedata),                  //          .writedata
		.rdclk_control_slave_write        (fifo_hps_to_fpga_out_csr_write),                      //          .write
		.rdclk_control_slave_readdata     (fifo_hps_to_fpga_out_csr_readdata),                   //          .readdata
		.wrclk_control_slave_address      (mm_interconnect_2_fifo_hps_to_fpga_in_csr_address),   //    in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_2_fifo_hps_to_fpga_in_csr_read),      //          .read
		.wrclk_control_slave_writedata    (mm_interconnect_2_fifo_hps_to_fpga_in_csr_writedata), //          .writedata
		.wrclk_control_slave_write        (mm_interconnect_2_fifo_hps_to_fpga_in_csr_write),     //          .write
		.wrclk_control_slave_readdata     (mm_interconnect_2_fifo_hps_to_fpga_in_csr_readdata)   //          .readdata
	);

	sys_vga_hex5_hex0 hex5_hex0 (
		.clk        (sys_sdram_pll_0_sys_clk_clk),               //                 clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_2_hex5_hex0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_hex5_hex0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_hex5_hex0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_hex5_hex0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_hex5_hex0_s1_readdata),   //                    .readdata
		.out_port   (hex5_0bus_export)                           // external_connection.export
	);

	sys_vga_new_sdram_controller_0 new_sdram_controller_0 (
		.clk            (sys_sdram_pll_0_sys_clk_clk),                               //   clk.clk
		.reset_n        (~rst_controller_003_reset_out_reset),                       // reset.reset_n
		.az_addr        (mm_interconnect_1_new_sdram_controller_0_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_1_new_sdram_controller_0_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_1_new_sdram_controller_0_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_1_new_sdram_controller_0_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_1_new_sdram_controller_0_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_1_new_sdram_controller_0_s1_write),        //      .write_n
		.za_data        (mm_interconnect_1_new_sdram_controller_0_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_1_new_sdram_controller_0_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_1_new_sdram_controller_0_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                                           //  wire.export
		.zs_ba          (sdram_wire_ba),                                             //      .export
		.zs_cas_n       (sdram_wire_cas_n),                                          //      .export
		.zs_cke         (sdram_wire_cke),                                            //      .export
		.zs_cs_n        (sdram_wire_cs_n),                                           //      .export
		.zs_dq          (sdram_wire_dq),                                             //      .export
		.zs_dqm         (sdram_wire_dqm),                                            //      .export
		.zs_ras_n       (sdram_wire_ras_n),                                          //      .export
		.zs_we_n        (sdram_wire_we_n)                                            //      .export
	);

	sys_vga_pll_0 pll_0 (
		.refclk   (sys_sdram_pll_0_sys_clk_clk),        //  refclk.clk
		.rst      (sys_sdram_pll_0_reset_source_reset), //   reset.reset
		.outclk_0 (pll_0_outclk0_clk),                  // outclk0.clk
		.locked   ()                                    //  locked.export
	);

	sys_vga_pll_1 pll_1 (
		.refclk   (sys_sdram_pll_0_sys_clk_clk),        //  refclk.clk
		.rst      (sys_sdram_pll_0_reset_source_reset), //   reset.reset
		.outclk_0 (clk_65_clk),                         // outclk0.clk
		.locked   ()                                    //  locked.export
	);

	sys_vga_pushbuttons pushbuttons (
		.clk        (sys_sdram_pll_0_sys_clk_clk),                 //                 clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_2_pushbuttons_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_pushbuttons_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_pushbuttons_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_pushbuttons_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_pushbuttons_s1_readdata),   //                    .readdata
		.in_port    (pushbutton_export),                           // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                     //                 irq.irq
	);

	sys_vga_ram ram (
		.clk         (sys_sdram_pll_0_sys_clk_clk),            //   clk1.clk
		.address     (mm_interconnect_1_ram_s1_address),       //     s1.address
		.clken       (mm_interconnect_1_ram_s1_clken),         //       .clken
		.chipselect  (mm_interconnect_1_ram_s1_chipselect),    //       .chipselect
		.write       (mm_interconnect_1_ram_s1_write),         //       .write
		.readdata    (mm_interconnect_1_ram_s1_readdata),      //       .readdata
		.writedata   (mm_interconnect_1_ram_s1_writedata),     //       .writedata
		.byteenable  (mm_interconnect_1_ram_s1_byteenable),    //       .byteenable
		.reset       (rst_controller_003_reset_out_reset),     // reset1.reset
		.reset_req   (rst_controller_003_reset_out_reset_req), //       .reset_req
		.address2    (ram_s2_address),                         //     s2.address
		.chipselect2 (ram_s2_chipselect),                      //       .chipselect
		.clken2      (ram_s2_clken),                           //       .clken
		.write2      (ram_s2_write),                           //       .write
		.readdata2   (ram_s2_readdata),                        //       .readdata
		.writedata2  (ram_s2_writedata),                       //       .writedata
		.byteenable2 (ram_s2_byteenable),                      //       .byteenable
		.clk2        (clock_bridge_0_in_clk_clk),              //   clk2.clk
		.reset2      (rst_controller_002_reset_out_reset),     // reset2.reset
		.reset_req2  (rst_controller_002_reset_out_reset_req), //       .reset_req
		.freeze      (1'b0)                                    // (terminated)
	);

	reg32_avalon_interface reg32_avalon_interface_0 (
		.clk        (sys_sdram_pll_0_sys_clk_clk),                                          //          clock.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                                  //          reset.reset_n
		.write      (mm_interconnect_2_reg32_avalon_interface_0_avalon_slave_0_write),      // avalon_slave_0.write
		.writedata  (mm_interconnect_2_reg32_avalon_interface_0_avalon_slave_0_writedata),  //               .writedata
		.read       (mm_interconnect_2_reg32_avalon_interface_0_avalon_slave_0_read),       //               .read
		.readdata   (mm_interconnect_2_reg32_avalon_interface_0_avalon_slave_0_readdata),   //               .readdata
		.byteenable (mm_interconnect_2_reg32_avalon_interface_0_avalon_slave_0_byteenable), //               .byteenable
		.chipselect (mm_interconnect_2_reg32_avalon_interface_0_avalon_slave_0_chipselect), //               .chipselect
		.Q_external (to_hex_to_led_readdata)                                                //    conduit_end.readdata
	);

	sys_vga_sys_sdram_pll_0 sys_sdram_pll_0 (
		.ref_clk_clk        (system_ref_clk_clk),                 //      ref_clk.clk
		.ref_reset_reset    (system_ref_reset_reset),             //    ref_reset.reset
		.sys_clk_clk        (sys_sdram_pll_0_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                      //    sdram_clk.clk
		.reset_source_reset (sys_sdram_pll_0_reset_source_reset)  // reset_source.reset
	);

	sys_vga_sysid_qsys_0 sysid_qsys_0 (
		.clock    (sys_sdram_pll_0_sys_clk_clk),                           //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_2_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_2_sysid_qsys_0_control_slave_address)   //              .address
	);

	sys_vga_system_console system_console (
		.clk            (sys_sdram_pll_0_sys_clk_clk),                                    //               clk.clk
		.rst_n          (~rst_controller_003_reset_out_reset),                            //             reset.reset_n
		.av_chipselect  (mm_interconnect_2_system_console_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_2_system_console_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_2_system_console_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_2_system_console_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_2_system_console_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_2_system_console_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_2_system_console_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                        //               irq.irq
	);

	sys_vga_mm_interconnect_0 mm_interconnect_0 (
		.Arm_A9_HPS_f2h_axi_slave_awid                                         (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awid),    //                                        Arm_A9_HPS_f2h_axi_slave.awid
		.Arm_A9_HPS_f2h_axi_slave_awaddr                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awaddr),  //                                                                .awaddr
		.Arm_A9_HPS_f2h_axi_slave_awlen                                        (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awlen),   //                                                                .awlen
		.Arm_A9_HPS_f2h_axi_slave_awsize                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awsize),  //                                                                .awsize
		.Arm_A9_HPS_f2h_axi_slave_awburst                                      (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awburst), //                                                                .awburst
		.Arm_A9_HPS_f2h_axi_slave_awlock                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awlock),  //                                                                .awlock
		.Arm_A9_HPS_f2h_axi_slave_awcache                                      (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awcache), //                                                                .awcache
		.Arm_A9_HPS_f2h_axi_slave_awprot                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awprot),  //                                                                .awprot
		.Arm_A9_HPS_f2h_axi_slave_awuser                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awuser),  //                                                                .awuser
		.Arm_A9_HPS_f2h_axi_slave_awvalid                                      (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awvalid), //                                                                .awvalid
		.Arm_A9_HPS_f2h_axi_slave_awready                                      (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_awready), //                                                                .awready
		.Arm_A9_HPS_f2h_axi_slave_wid                                          (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wid),     //                                                                .wid
		.Arm_A9_HPS_f2h_axi_slave_wdata                                        (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wdata),   //                                                                .wdata
		.Arm_A9_HPS_f2h_axi_slave_wstrb                                        (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wstrb),   //                                                                .wstrb
		.Arm_A9_HPS_f2h_axi_slave_wlast                                        (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wlast),   //                                                                .wlast
		.Arm_A9_HPS_f2h_axi_slave_wvalid                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wvalid),  //                                                                .wvalid
		.Arm_A9_HPS_f2h_axi_slave_wready                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_wready),  //                                                                .wready
		.Arm_A9_HPS_f2h_axi_slave_bid                                          (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bid),     //                                                                .bid
		.Arm_A9_HPS_f2h_axi_slave_bresp                                        (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bresp),   //                                                                .bresp
		.Arm_A9_HPS_f2h_axi_slave_bvalid                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bvalid),  //                                                                .bvalid
		.Arm_A9_HPS_f2h_axi_slave_bready                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_bready),  //                                                                .bready
		.Arm_A9_HPS_f2h_axi_slave_arid                                         (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arid),    //                                                                .arid
		.Arm_A9_HPS_f2h_axi_slave_araddr                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_araddr),  //                                                                .araddr
		.Arm_A9_HPS_f2h_axi_slave_arlen                                        (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arlen),   //                                                                .arlen
		.Arm_A9_HPS_f2h_axi_slave_arsize                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arsize),  //                                                                .arsize
		.Arm_A9_HPS_f2h_axi_slave_arburst                                      (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arburst), //                                                                .arburst
		.Arm_A9_HPS_f2h_axi_slave_arlock                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arlock),  //                                                                .arlock
		.Arm_A9_HPS_f2h_axi_slave_arcache                                      (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arcache), //                                                                .arcache
		.Arm_A9_HPS_f2h_axi_slave_arprot                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arprot),  //                                                                .arprot
		.Arm_A9_HPS_f2h_axi_slave_aruser                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_aruser),  //                                                                .aruser
		.Arm_A9_HPS_f2h_axi_slave_arvalid                                      (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arvalid), //                                                                .arvalid
		.Arm_A9_HPS_f2h_axi_slave_arready                                      (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_arready), //                                                                .arready
		.Arm_A9_HPS_f2h_axi_slave_rid                                          (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rid),     //                                                                .rid
		.Arm_A9_HPS_f2h_axi_slave_rdata                                        (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rdata),   //                                                                .rdata
		.Arm_A9_HPS_f2h_axi_slave_rresp                                        (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rresp),   //                                                                .rresp
		.Arm_A9_HPS_f2h_axi_slave_rlast                                        (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rlast),   //                                                                .rlast
		.Arm_A9_HPS_f2h_axi_slave_rvalid                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rvalid),  //                                                                .rvalid
		.Arm_A9_HPS_f2h_axi_slave_rready                                       (mm_interconnect_0_arm_a9_hps_f2h_axi_slave_rready),  //                                                                .rready
		.sys_sdram_pll_0_sys_clk_clk                                           (sys_sdram_pll_0_sys_clk_clk),                        //                                         sys_sdram_pll_0_sys_clk.clk
		.alt_vip_vfr_0_clock_master_reset_reset_bridge_in_reset_reset          (rst_controller_001_reset_out_reset),                 //          alt_vip_vfr_0_clock_master_reset_reset_bridge_in_reset.reset
		.Arm_A9_HPS_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset (rst_controller_004_reset_out_reset),                 // Arm_A9_HPS_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset.reset
		.alt_vip_vfr_0_avalon_master_address                                   (alt_vip_vfr_0_avalon_master_address),                //                                     alt_vip_vfr_0_avalon_master.address
		.alt_vip_vfr_0_avalon_master_waitrequest                               (alt_vip_vfr_0_avalon_master_waitrequest),            //                                                                .waitrequest
		.alt_vip_vfr_0_avalon_master_burstcount                                (alt_vip_vfr_0_avalon_master_burstcount),             //                                                                .burstcount
		.alt_vip_vfr_0_avalon_master_read                                      (alt_vip_vfr_0_avalon_master_read),                   //                                                                .read
		.alt_vip_vfr_0_avalon_master_readdata                                  (alt_vip_vfr_0_avalon_master_readdata),               //                                                                .readdata
		.alt_vip_vfr_0_avalon_master_readdatavalid                             (alt_vip_vfr_0_avalon_master_readdatavalid)           //                                                                .readdatavalid
	);

	sys_vga_mm_interconnect_1 mm_interconnect_1 (
		.Arm_A9_HPS_h2f_axi_master_awid                                        (arm_a9_hps_h2f_axi_master_awid),                            //                                       Arm_A9_HPS_h2f_axi_master.awid
		.Arm_A9_HPS_h2f_axi_master_awaddr                                      (arm_a9_hps_h2f_axi_master_awaddr),                          //                                                                .awaddr
		.Arm_A9_HPS_h2f_axi_master_awlen                                       (arm_a9_hps_h2f_axi_master_awlen),                           //                                                                .awlen
		.Arm_A9_HPS_h2f_axi_master_awsize                                      (arm_a9_hps_h2f_axi_master_awsize),                          //                                                                .awsize
		.Arm_A9_HPS_h2f_axi_master_awburst                                     (arm_a9_hps_h2f_axi_master_awburst),                         //                                                                .awburst
		.Arm_A9_HPS_h2f_axi_master_awlock                                      (arm_a9_hps_h2f_axi_master_awlock),                          //                                                                .awlock
		.Arm_A9_HPS_h2f_axi_master_awcache                                     (arm_a9_hps_h2f_axi_master_awcache),                         //                                                                .awcache
		.Arm_A9_HPS_h2f_axi_master_awprot                                      (arm_a9_hps_h2f_axi_master_awprot),                          //                                                                .awprot
		.Arm_A9_HPS_h2f_axi_master_awvalid                                     (arm_a9_hps_h2f_axi_master_awvalid),                         //                                                                .awvalid
		.Arm_A9_HPS_h2f_axi_master_awready                                     (arm_a9_hps_h2f_axi_master_awready),                         //                                                                .awready
		.Arm_A9_HPS_h2f_axi_master_wid                                         (arm_a9_hps_h2f_axi_master_wid),                             //                                                                .wid
		.Arm_A9_HPS_h2f_axi_master_wdata                                       (arm_a9_hps_h2f_axi_master_wdata),                           //                                                                .wdata
		.Arm_A9_HPS_h2f_axi_master_wstrb                                       (arm_a9_hps_h2f_axi_master_wstrb),                           //                                                                .wstrb
		.Arm_A9_HPS_h2f_axi_master_wlast                                       (arm_a9_hps_h2f_axi_master_wlast),                           //                                                                .wlast
		.Arm_A9_HPS_h2f_axi_master_wvalid                                      (arm_a9_hps_h2f_axi_master_wvalid),                          //                                                                .wvalid
		.Arm_A9_HPS_h2f_axi_master_wready                                      (arm_a9_hps_h2f_axi_master_wready),                          //                                                                .wready
		.Arm_A9_HPS_h2f_axi_master_bid                                         (arm_a9_hps_h2f_axi_master_bid),                             //                                                                .bid
		.Arm_A9_HPS_h2f_axi_master_bresp                                       (arm_a9_hps_h2f_axi_master_bresp),                           //                                                                .bresp
		.Arm_A9_HPS_h2f_axi_master_bvalid                                      (arm_a9_hps_h2f_axi_master_bvalid),                          //                                                                .bvalid
		.Arm_A9_HPS_h2f_axi_master_bready                                      (arm_a9_hps_h2f_axi_master_bready),                          //                                                                .bready
		.Arm_A9_HPS_h2f_axi_master_arid                                        (arm_a9_hps_h2f_axi_master_arid),                            //                                                                .arid
		.Arm_A9_HPS_h2f_axi_master_araddr                                      (arm_a9_hps_h2f_axi_master_araddr),                          //                                                                .araddr
		.Arm_A9_HPS_h2f_axi_master_arlen                                       (arm_a9_hps_h2f_axi_master_arlen),                           //                                                                .arlen
		.Arm_A9_HPS_h2f_axi_master_arsize                                      (arm_a9_hps_h2f_axi_master_arsize),                          //                                                                .arsize
		.Arm_A9_HPS_h2f_axi_master_arburst                                     (arm_a9_hps_h2f_axi_master_arburst),                         //                                                                .arburst
		.Arm_A9_HPS_h2f_axi_master_arlock                                      (arm_a9_hps_h2f_axi_master_arlock),                          //                                                                .arlock
		.Arm_A9_HPS_h2f_axi_master_arcache                                     (arm_a9_hps_h2f_axi_master_arcache),                         //                                                                .arcache
		.Arm_A9_HPS_h2f_axi_master_arprot                                      (arm_a9_hps_h2f_axi_master_arprot),                          //                                                                .arprot
		.Arm_A9_HPS_h2f_axi_master_arvalid                                     (arm_a9_hps_h2f_axi_master_arvalid),                         //                                                                .arvalid
		.Arm_A9_HPS_h2f_axi_master_arready                                     (arm_a9_hps_h2f_axi_master_arready),                         //                                                                .arready
		.Arm_A9_HPS_h2f_axi_master_rid                                         (arm_a9_hps_h2f_axi_master_rid),                             //                                                                .rid
		.Arm_A9_HPS_h2f_axi_master_rdata                                       (arm_a9_hps_h2f_axi_master_rdata),                           //                                                                .rdata
		.Arm_A9_HPS_h2f_axi_master_rresp                                       (arm_a9_hps_h2f_axi_master_rresp),                           //                                                                .rresp
		.Arm_A9_HPS_h2f_axi_master_rlast                                       (arm_a9_hps_h2f_axi_master_rlast),                           //                                                                .rlast
		.Arm_A9_HPS_h2f_axi_master_rvalid                                      (arm_a9_hps_h2f_axi_master_rvalid),                          //                                                                .rvalid
		.Arm_A9_HPS_h2f_axi_master_rready                                      (arm_a9_hps_h2f_axi_master_rready),                          //                                                                .rready
		.sys_sdram_pll_0_sys_clk_clk                                           (sys_sdram_pll_0_sys_clk_clk),                               //                                         sys_sdram_pll_0_sys_clk.clk
		.Arm_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_004_reset_out_reset),                        // Arm_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.fifo_hps_to_fpga_reset_in_reset_bridge_in_reset_reset                 (rst_controller_003_reset_out_reset),                        //                 fifo_hps_to_fpga_reset_in_reset_bridge_in_reset.reset
		.fifo_fpga_to_hps_out_read                                             (mm_interconnect_1_fifo_fpga_to_hps_out_read),               //                                            fifo_fpga_to_hps_out.read
		.fifo_fpga_to_hps_out_readdata                                         (mm_interconnect_1_fifo_fpga_to_hps_out_readdata),           //                                                                .readdata
		.fifo_fpga_to_hps_out_waitrequest                                      (mm_interconnect_1_fifo_fpga_to_hps_out_waitrequest),        //                                                                .waitrequest
		.fifo_hps_to_fpga_in_write                                             (mm_interconnect_1_fifo_hps_to_fpga_in_write),               //                                             fifo_hps_to_fpga_in.write
		.fifo_hps_to_fpga_in_writedata                                         (mm_interconnect_1_fifo_hps_to_fpga_in_writedata),           //                                                                .writedata
		.fifo_hps_to_fpga_in_waitrequest                                       (mm_interconnect_1_fifo_hps_to_fpga_in_waitrequest),         //                                                                .waitrequest
		.new_sdram_controller_0_s1_address                                     (mm_interconnect_1_new_sdram_controller_0_s1_address),       //                                       new_sdram_controller_0_s1.address
		.new_sdram_controller_0_s1_write                                       (mm_interconnect_1_new_sdram_controller_0_s1_write),         //                                                                .write
		.new_sdram_controller_0_s1_read                                        (mm_interconnect_1_new_sdram_controller_0_s1_read),          //                                                                .read
		.new_sdram_controller_0_s1_readdata                                    (mm_interconnect_1_new_sdram_controller_0_s1_readdata),      //                                                                .readdata
		.new_sdram_controller_0_s1_writedata                                   (mm_interconnect_1_new_sdram_controller_0_s1_writedata),     //                                                                .writedata
		.new_sdram_controller_0_s1_byteenable                                  (mm_interconnect_1_new_sdram_controller_0_s1_byteenable),    //                                                                .byteenable
		.new_sdram_controller_0_s1_readdatavalid                               (mm_interconnect_1_new_sdram_controller_0_s1_readdatavalid), //                                                                .readdatavalid
		.new_sdram_controller_0_s1_waitrequest                                 (mm_interconnect_1_new_sdram_controller_0_s1_waitrequest),   //                                                                .waitrequest
		.new_sdram_controller_0_s1_chipselect                                  (mm_interconnect_1_new_sdram_controller_0_s1_chipselect),    //                                                                .chipselect
		.ram_s1_address                                                        (mm_interconnect_1_ram_s1_address),                          //                                                          ram_s1.address
		.ram_s1_write                                                          (mm_interconnect_1_ram_s1_write),                            //                                                                .write
		.ram_s1_readdata                                                       (mm_interconnect_1_ram_s1_readdata),                         //                                                                .readdata
		.ram_s1_writedata                                                      (mm_interconnect_1_ram_s1_writedata),                        //                                                                .writedata
		.ram_s1_byteenable                                                     (mm_interconnect_1_ram_s1_byteenable),                       //                                                                .byteenable
		.ram_s1_chipselect                                                     (mm_interconnect_1_ram_s1_chipselect),                       //                                                                .chipselect
		.ram_s1_clken                                                          (mm_interconnect_1_ram_s1_clken)                             //                                                                .clken
	);

	sys_vga_mm_interconnect_2 mm_interconnect_2 (
		.Arm_A9_HPS_h2f_lw_axi_master_awid                                        (arm_a9_hps_h2f_lw_axi_master_awid),                                    //                                       Arm_A9_HPS_h2f_lw_axi_master.awid
		.Arm_A9_HPS_h2f_lw_axi_master_awaddr                                      (arm_a9_hps_h2f_lw_axi_master_awaddr),                                  //                                                                   .awaddr
		.Arm_A9_HPS_h2f_lw_axi_master_awlen                                       (arm_a9_hps_h2f_lw_axi_master_awlen),                                   //                                                                   .awlen
		.Arm_A9_HPS_h2f_lw_axi_master_awsize                                      (arm_a9_hps_h2f_lw_axi_master_awsize),                                  //                                                                   .awsize
		.Arm_A9_HPS_h2f_lw_axi_master_awburst                                     (arm_a9_hps_h2f_lw_axi_master_awburst),                                 //                                                                   .awburst
		.Arm_A9_HPS_h2f_lw_axi_master_awlock                                      (arm_a9_hps_h2f_lw_axi_master_awlock),                                  //                                                                   .awlock
		.Arm_A9_HPS_h2f_lw_axi_master_awcache                                     (arm_a9_hps_h2f_lw_axi_master_awcache),                                 //                                                                   .awcache
		.Arm_A9_HPS_h2f_lw_axi_master_awprot                                      (arm_a9_hps_h2f_lw_axi_master_awprot),                                  //                                                                   .awprot
		.Arm_A9_HPS_h2f_lw_axi_master_awvalid                                     (arm_a9_hps_h2f_lw_axi_master_awvalid),                                 //                                                                   .awvalid
		.Arm_A9_HPS_h2f_lw_axi_master_awready                                     (arm_a9_hps_h2f_lw_axi_master_awready),                                 //                                                                   .awready
		.Arm_A9_HPS_h2f_lw_axi_master_wid                                         (arm_a9_hps_h2f_lw_axi_master_wid),                                     //                                                                   .wid
		.Arm_A9_HPS_h2f_lw_axi_master_wdata                                       (arm_a9_hps_h2f_lw_axi_master_wdata),                                   //                                                                   .wdata
		.Arm_A9_HPS_h2f_lw_axi_master_wstrb                                       (arm_a9_hps_h2f_lw_axi_master_wstrb),                                   //                                                                   .wstrb
		.Arm_A9_HPS_h2f_lw_axi_master_wlast                                       (arm_a9_hps_h2f_lw_axi_master_wlast),                                   //                                                                   .wlast
		.Arm_A9_HPS_h2f_lw_axi_master_wvalid                                      (arm_a9_hps_h2f_lw_axi_master_wvalid),                                  //                                                                   .wvalid
		.Arm_A9_HPS_h2f_lw_axi_master_wready                                      (arm_a9_hps_h2f_lw_axi_master_wready),                                  //                                                                   .wready
		.Arm_A9_HPS_h2f_lw_axi_master_bid                                         (arm_a9_hps_h2f_lw_axi_master_bid),                                     //                                                                   .bid
		.Arm_A9_HPS_h2f_lw_axi_master_bresp                                       (arm_a9_hps_h2f_lw_axi_master_bresp),                                   //                                                                   .bresp
		.Arm_A9_HPS_h2f_lw_axi_master_bvalid                                      (arm_a9_hps_h2f_lw_axi_master_bvalid),                                  //                                                                   .bvalid
		.Arm_A9_HPS_h2f_lw_axi_master_bready                                      (arm_a9_hps_h2f_lw_axi_master_bready),                                  //                                                                   .bready
		.Arm_A9_HPS_h2f_lw_axi_master_arid                                        (arm_a9_hps_h2f_lw_axi_master_arid),                                    //                                                                   .arid
		.Arm_A9_HPS_h2f_lw_axi_master_araddr                                      (arm_a9_hps_h2f_lw_axi_master_araddr),                                  //                                                                   .araddr
		.Arm_A9_HPS_h2f_lw_axi_master_arlen                                       (arm_a9_hps_h2f_lw_axi_master_arlen),                                   //                                                                   .arlen
		.Arm_A9_HPS_h2f_lw_axi_master_arsize                                      (arm_a9_hps_h2f_lw_axi_master_arsize),                                  //                                                                   .arsize
		.Arm_A9_HPS_h2f_lw_axi_master_arburst                                     (arm_a9_hps_h2f_lw_axi_master_arburst),                                 //                                                                   .arburst
		.Arm_A9_HPS_h2f_lw_axi_master_arlock                                      (arm_a9_hps_h2f_lw_axi_master_arlock),                                  //                                                                   .arlock
		.Arm_A9_HPS_h2f_lw_axi_master_arcache                                     (arm_a9_hps_h2f_lw_axi_master_arcache),                                 //                                                                   .arcache
		.Arm_A9_HPS_h2f_lw_axi_master_arprot                                      (arm_a9_hps_h2f_lw_axi_master_arprot),                                  //                                                                   .arprot
		.Arm_A9_HPS_h2f_lw_axi_master_arvalid                                     (arm_a9_hps_h2f_lw_axi_master_arvalid),                                 //                                                                   .arvalid
		.Arm_A9_HPS_h2f_lw_axi_master_arready                                     (arm_a9_hps_h2f_lw_axi_master_arready),                                 //                                                                   .arready
		.Arm_A9_HPS_h2f_lw_axi_master_rid                                         (arm_a9_hps_h2f_lw_axi_master_rid),                                     //                                                                   .rid
		.Arm_A9_HPS_h2f_lw_axi_master_rdata                                       (arm_a9_hps_h2f_lw_axi_master_rdata),                                   //                                                                   .rdata
		.Arm_A9_HPS_h2f_lw_axi_master_rresp                                       (arm_a9_hps_h2f_lw_axi_master_rresp),                                   //                                                                   .rresp
		.Arm_A9_HPS_h2f_lw_axi_master_rlast                                       (arm_a9_hps_h2f_lw_axi_master_rlast),                                   //                                                                   .rlast
		.Arm_A9_HPS_h2f_lw_axi_master_rvalid                                      (arm_a9_hps_h2f_lw_axi_master_rvalid),                                  //                                                                   .rvalid
		.Arm_A9_HPS_h2f_lw_axi_master_rready                                      (arm_a9_hps_h2f_lw_axi_master_rready),                                  //                                                                   .rready
		.pll_0_outclk0_clk                                                        (pll_0_outclk0_clk),                                                    //                                                      pll_0_outclk0.clk
		.sys_sdram_pll_0_sys_clk_clk                                              (sys_sdram_pll_0_sys_clk_clk),                                          //                                            sys_sdram_pll_0_sys_clk.clk
		.alt_vip_vfr_0_clock_reset_reset_reset_bridge_in_reset_reset              (rst_controller_reset_out_reset),                                       //              alt_vip_vfr_0_clock_reset_reset_reset_bridge_in_reset.reset
		.Arm_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_004_reset_out_reset),                                   // Arm_A9_HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.sysid_qsys_0_reset_reset_bridge_in_reset_reset                           (rst_controller_001_reset_out_reset),                                   //                           sysid_qsys_0_reset_reset_bridge_in_reset.reset
		.system_console_reset_reset_bridge_in_reset_reset                         (rst_controller_003_reset_out_reset),                                   //                         system_console_reset_reset_bridge_in_reset.reset
		.alt_vip_vfr_0_avalon_slave_address                                       (mm_interconnect_2_alt_vip_vfr_0_avalon_slave_address),                 //                                         alt_vip_vfr_0_avalon_slave.address
		.alt_vip_vfr_0_avalon_slave_write                                         (mm_interconnect_2_alt_vip_vfr_0_avalon_slave_write),                   //                                                                   .write
		.alt_vip_vfr_0_avalon_slave_read                                          (mm_interconnect_2_alt_vip_vfr_0_avalon_slave_read),                    //                                                                   .read
		.alt_vip_vfr_0_avalon_slave_readdata                                      (mm_interconnect_2_alt_vip_vfr_0_avalon_slave_readdata),                //                                                                   .readdata
		.alt_vip_vfr_0_avalon_slave_writedata                                     (mm_interconnect_2_alt_vip_vfr_0_avalon_slave_writedata),               //                                                                   .writedata
		.fifo_fpga_to_hps_out_csr_address                                         (mm_interconnect_2_fifo_fpga_to_hps_out_csr_address),                   //                                           fifo_fpga_to_hps_out_csr.address
		.fifo_fpga_to_hps_out_csr_write                                           (mm_interconnect_2_fifo_fpga_to_hps_out_csr_write),                     //                                                                   .write
		.fifo_fpga_to_hps_out_csr_read                                            (mm_interconnect_2_fifo_fpga_to_hps_out_csr_read),                      //                                                                   .read
		.fifo_fpga_to_hps_out_csr_readdata                                        (mm_interconnect_2_fifo_fpga_to_hps_out_csr_readdata),                  //                                                                   .readdata
		.fifo_fpga_to_hps_out_csr_writedata                                       (mm_interconnect_2_fifo_fpga_to_hps_out_csr_writedata),                 //                                                                   .writedata
		.fifo_hps_to_fpga_in_csr_address                                          (mm_interconnect_2_fifo_hps_to_fpga_in_csr_address),                    //                                            fifo_hps_to_fpga_in_csr.address
		.fifo_hps_to_fpga_in_csr_write                                            (mm_interconnect_2_fifo_hps_to_fpga_in_csr_write),                      //                                                                   .write
		.fifo_hps_to_fpga_in_csr_read                                             (mm_interconnect_2_fifo_hps_to_fpga_in_csr_read),                       //                                                                   .read
		.fifo_hps_to_fpga_in_csr_readdata                                         (mm_interconnect_2_fifo_hps_to_fpga_in_csr_readdata),                   //                                                                   .readdata
		.fifo_hps_to_fpga_in_csr_writedata                                        (mm_interconnect_2_fifo_hps_to_fpga_in_csr_writedata),                  //                                                                   .writedata
		.hex5_hex0_s1_address                                                     (mm_interconnect_2_hex5_hex0_s1_address),                               //                                                       hex5_hex0_s1.address
		.hex5_hex0_s1_write                                                       (mm_interconnect_2_hex5_hex0_s1_write),                                 //                                                                   .write
		.hex5_hex0_s1_readdata                                                    (mm_interconnect_2_hex5_hex0_s1_readdata),                              //                                                                   .readdata
		.hex5_hex0_s1_writedata                                                   (mm_interconnect_2_hex5_hex0_s1_writedata),                             //                                                                   .writedata
		.hex5_hex0_s1_chipselect                                                  (mm_interconnect_2_hex5_hex0_s1_chipselect),                            //                                                                   .chipselect
		.pushbuttons_s1_address                                                   (mm_interconnect_2_pushbuttons_s1_address),                             //                                                     pushbuttons_s1.address
		.pushbuttons_s1_write                                                     (mm_interconnect_2_pushbuttons_s1_write),                               //                                                                   .write
		.pushbuttons_s1_readdata                                                  (mm_interconnect_2_pushbuttons_s1_readdata),                            //                                                                   .readdata
		.pushbuttons_s1_writedata                                                 (mm_interconnect_2_pushbuttons_s1_writedata),                           //                                                                   .writedata
		.pushbuttons_s1_chipselect                                                (mm_interconnect_2_pushbuttons_s1_chipselect),                          //                                                                   .chipselect
		.reg32_avalon_interface_0_avalon_slave_0_write                            (mm_interconnect_2_reg32_avalon_interface_0_avalon_slave_0_write),      //                            reg32_avalon_interface_0_avalon_slave_0.write
		.reg32_avalon_interface_0_avalon_slave_0_read                             (mm_interconnect_2_reg32_avalon_interface_0_avalon_slave_0_read),       //                                                                   .read
		.reg32_avalon_interface_0_avalon_slave_0_readdata                         (mm_interconnect_2_reg32_avalon_interface_0_avalon_slave_0_readdata),   //                                                                   .readdata
		.reg32_avalon_interface_0_avalon_slave_0_writedata                        (mm_interconnect_2_reg32_avalon_interface_0_avalon_slave_0_writedata),  //                                                                   .writedata
		.reg32_avalon_interface_0_avalon_slave_0_byteenable                       (mm_interconnect_2_reg32_avalon_interface_0_avalon_slave_0_byteenable), //                                                                   .byteenable
		.reg32_avalon_interface_0_avalon_slave_0_chipselect                       (mm_interconnect_2_reg32_avalon_interface_0_avalon_slave_0_chipselect), //                                                                   .chipselect
		.sysid_qsys_0_control_slave_address                                       (mm_interconnect_2_sysid_qsys_0_control_slave_address),                 //                                         sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                                      (mm_interconnect_2_sysid_qsys_0_control_slave_readdata),                //                                                                   .readdata
		.system_console_avalon_jtag_slave_address                                 (mm_interconnect_2_system_console_avalon_jtag_slave_address),           //                                   system_console_avalon_jtag_slave.address
		.system_console_avalon_jtag_slave_write                                   (mm_interconnect_2_system_console_avalon_jtag_slave_write),             //                                                                   .write
		.system_console_avalon_jtag_slave_read                                    (mm_interconnect_2_system_console_avalon_jtag_slave_read),              //                                                                   .read
		.system_console_avalon_jtag_slave_readdata                                (mm_interconnect_2_system_console_avalon_jtag_slave_readdata),          //                                                                   .readdata
		.system_console_avalon_jtag_slave_writedata                               (mm_interconnect_2_system_console_avalon_jtag_slave_writedata),         //                                                                   .writedata
		.system_console_avalon_jtag_slave_waitrequest                             (mm_interconnect_2_system_console_avalon_jtag_slave_waitrequest),       //                                                                   .waitrequest
		.system_console_avalon_jtag_slave_chipselect                              (mm_interconnect_2_system_console_avalon_jtag_slave_chipselect)         //                                                                   .chipselect
	);

	sys_vga_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq), // receiver1.irq
		.sender_irq    (arm_a9_hps_f2h_irq0_irq)   //    sender.irq
	);

	sys_vga_irq_mapper_001 irq_mapper_001 (
		.clk        (),                        //       clk.clk
		.reset      (),                        // clk_reset.reset
		.sender_irq (arm_a9_hps_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (sys_sdram_pll_0_reset_source_reset), // reset_in0.reset
		.clk            (pll_0_outclk0_clk),                  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (sys_sdram_pll_0_reset_source_reset), // reset_in0.reset
		.clk            (sys_sdram_pll_0_sys_clk_clk),        //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),            // reset_in0.reset
		.reset_in1      (sys_sdram_pll_0_reset_source_reset),     // reset_in1.reset
		.clk            (clock_bridge_0_in_clk_clk),              //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),            // reset_in0.reset
		.reset_in1      (sys_sdram_pll_0_reset_source_reset),     // reset_in1.reset
		.clk            (sys_sdram_pll_0_sys_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_003_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.clk            (sys_sdram_pll_0_sys_clk_clk),        //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
